
module Rom(output reg[11:0] out, input[10:0] address, input clk);
 
always @(posedge clk)
 begin	

	  case(address)	
270 : out <= 12'b001000100010;
271 : out <= 12'b001000100001;
272 : out <= 12'b001000100000;
273 : out <= 12'b001000011001;
274 : out <= 12'b001000011000;
275 : out <= 12'b001000011000;
276 : out <= 12'b001000010111;
277 : out <= 12'b001000010110;
278 : out <= 12'b001000010101;
279 : out <= 12'b001000010101;
280 : out <= 12'b001000010100;
281 : out <= 12'b001000010011;
282 : out <= 12'b001000010010;
283 : out <= 12'b001000010010;
284 : out <= 12'b001000010001;
285 : out <= 12'b001000010000;
286 : out <= 12'b001000001001;
287 : out <= 12'b001000001001;
288 : out <= 12'b001000001000;
289 : out <= 12'b001000000111;
290 : out <= 12'b001000000110;
291 : out <= 12'b001000000110;
292 : out <= 12'b001000000101;
293 : out <= 12'b001000000100;
294 : out <= 12'b001000000100;
295 : out <= 12'b001000000011;
296 : out <= 12'b001000000010;
297 : out <= 12'b001000000010;
298 : out <= 12'b001000000001;
299 : out <= 12'b001000000000;
300 : out <= 12'b001000000000;
301 : out <= 12'b000110011001;
302 : out <= 12'b000110011000;
303 : out <= 12'b000110011000;
304 : out <= 12'b000110010111;
305 : out <= 12'b000110010110;
306 : out <= 12'b000110010110;
307 : out <= 12'b000110010101;
308 : out <= 12'b000110010100;
309 : out <= 12'b000110010100;
310 : out <= 12'b000110010011;
311 : out <= 12'b000110010010;
312 : out <= 12'b000110010010;
313 : out <= 12'b000110010001;
314 : out <= 12'b000110010001;
315 : out <= 12'b000110010000;
316 : out <= 12'b000110001001;
317 : out <= 12'b000110001001;
318 : out <= 12'b000110001000;
319 : out <= 12'b000110001000;
320 : out <= 12'b000110000111;
321 : out <= 12'b000110000110;
322 : out <= 12'b000110000110;
323 : out <= 12'b000110000101;
324 : out <= 12'b000110000101;
325 : out <= 12'b000110000100;
326 : out <= 12'b000110000100;
327 : out <= 12'b000110000011;
328 : out <= 12'b000110000010;
329 : out <= 12'b000110000010;
330 : out <= 12'b000110000001;
331 : out <= 12'b000110000001;
332 : out <= 12'b000110000000;
333 : out <= 12'b000110000000;
334 : out <= 12'b000101111001;
335 : out <= 12'b000101111001;
336 : out <= 12'b000101111000;
337 : out <= 12'b000101111000;
338 : out <= 12'b000101110111;
339 : out <= 12'b000101110110;
340 : out <= 12'b000101110110;
341 : out <= 12'b000101110101;
342 : out <= 12'b000101110101;
343 : out <= 12'b000101110100;
344 : out <= 12'b000101110100;
345 : out <= 12'b000101110011;
346 : out <= 12'b000101110011;
347 : out <= 12'b000101110010;
348 : out <= 12'b000101110010;
349 : out <= 12'b000101110001;
350 : out <= 12'b000101110001;
351 : out <= 12'b000101110000;
352 : out <= 12'b000101110000;
353 : out <= 12'b000101101001;
354 : out <= 12'b000101101001;
355 : out <= 12'b000101101001;
356 : out <= 12'b000101101000;
357 : out <= 12'b000101101000;
358 : out <= 12'b000101100111;
359 : out <= 12'b000101100111;
360 : out <= 12'b000101100110;
361 : out <= 12'b000101100110;
362 : out <= 12'b000101100101;
363 : out <= 12'b000101100101;
364 : out <= 12'b000101100100;
365 : out <= 12'b000101100100;
366 : out <= 12'b000101100011;
367 : out <= 12'b000101100011;
368 : out <= 12'b000101100011;
369 : out <= 12'b000101100010;
370 : out <= 12'b000101100010;
371 : out <= 12'b000101100001;
372 : out <= 12'b000101100001;
373 : out <= 12'b000101100000;
374 : out <= 12'b000101100000;
375 : out <= 12'b000101100000;
376 : out <= 12'b000101011001;
377 : out <= 12'b000101011001;
378 : out <= 12'b000101011000;
379 : out <= 12'b000101011000;
380 : out <= 12'b000101010111;
381 : out <= 12'b000101010111;
382 : out <= 12'b000101010111;
383 : out <= 12'b000101010110;
384 : out <= 12'b000101010110;
385 : out <= 12'b000101010101;
386 : out <= 12'b000101010101;
387 : out <= 12'b000101010101;
388 : out <= 12'b000101010100;
389 : out <= 12'b000101010100;
390 : out <= 12'b000101010011;
391 : out <= 12'b000101010011;
392 : out <= 12'b000101010011;
393 : out <= 12'b000101010010;
394 : out <= 12'b000101010010;
395 : out <= 12'b000101010001;
396 : out <= 12'b000101010001;
397 : out <= 12'b000101010001;
398 : out <= 12'b000101010000;
399 : out <= 12'b000101010000;
400 : out <= 12'b000101010000;
401 : out <= 12'b000101001001;
402 : out <= 12'b000101001001;
403 : out <= 12'b000101001000;
404 : out <= 12'b000101001000;
405 : out <= 12'b000101001000;
406 : out <= 12'b000101000111;
407 : out <= 12'b000101000111;
408 : out <= 12'b000101000111;
409 : out <= 12'b000101000110;
410 : out <= 12'b000101000110;
411 : out <= 12'b000101000101;
412 : out <= 12'b000101000101;
413 : out <= 12'b000101000101;
414 : out <= 12'b000101000100;
415 : out <= 12'b000101000100;
416 : out <= 12'b000101000100;
417 : out <= 12'b000101000011;
418 : out <= 12'b000101000011;
419 : out <= 12'b000101000011;
420 : out <= 12'b000101000010;
421 : out <= 12'b000101000010;
422 : out <= 12'b000101000010;
423 : out <= 12'b000101000001;
424 : out <= 12'b000101000001;
425 : out <= 12'b000101000001;
426 : out <= 12'b000101000000;
427 : out <= 12'b000101000000;
428 : out <= 12'b000101000000;
429 : out <= 12'b000100111001;
430 : out <= 12'b000100111001;
431 : out <= 12'b000100111001;
432 : out <= 12'b000100111000;
433 : out <= 12'b000100111000;
434 : out <= 12'b000100111000;
435 : out <= 12'b000100110111;
436 : out <= 12'b000100110111;
437 : out <= 12'b000100110111;
438 : out <= 12'b000100110110;
439 : out <= 12'b000100110110;
440 : out <= 12'b000100110110;
441 : out <= 12'b000100110110;
442 : out <= 12'b000100110101;
443 : out <= 12'b000100110101;
444 : out <= 12'b000100110101;
445 : out <= 12'b000100110100;
446 : out <= 12'b000100110100;
447 : out <= 12'b000100110100;
448 : out <= 12'b000100110011;
449 : out <= 12'b000100110011;
450 : out <= 12'b000100110011;
451 : out <= 12'b000100110011;
452 : out <= 12'b000100110010;
453 : out <= 12'b000100110010;
454 : out <= 12'b000100110010;
455 : out <= 12'b000100110001;
456 : out <= 12'b000100110001;
457 : out <= 12'b000100110001;
458 : out <= 12'b000100110001;
459 : out <= 12'b000100110000;
460 : out <= 12'b000100110000;
461 : out <= 12'b000100110000;
462 : out <= 12'b000100101001;
463 : out <= 12'b000100101001;
464 : out <= 12'b000100101001;
465 : out <= 12'b000100101001;
466 : out <= 12'b000100101000;
467 : out <= 12'b000100101000;
468 : out <= 12'b000100101000;
469 : out <= 12'b000100100111;
470 : out <= 12'b000100100111;
471 : out <= 12'b000100100111;
472 : out <= 12'b000100100111;
473 : out <= 12'b000100100110;
474 : out <= 12'b000100100110;
475 : out <= 12'b000100100110;
476 : out <= 12'b000100100110;
477 : out <= 12'b000100100101;
478 : out <= 12'b000100100101;
479 : out <= 12'b000100100101;
480 : out <= 12'b000100100101;
481 : out <= 12'b000100100100;
482 : out <= 12'b000100100100;
483 : out <= 12'b000100100100;
484 : out <= 12'b000100100011;
485 : out <= 12'b000100100011;
486 : out <= 12'b000100100011;
487 : out <= 12'b000100100011;
488 : out <= 12'b000100100010;
489 : out <= 12'b000100100010;
490 : out <= 12'b000100100010;
491 : out <= 12'b000100100010;
492 : out <= 12'b000100100001;
493 : out <= 12'b000100100001;
494 : out <= 12'b000100100001;
495 : out <= 12'b000100100001;
496 : out <= 12'b000100100000;
497 : out <= 12'b000100100000;
498 : out <= 12'b000100100000;
499 : out <= 12'b000100100000;
500 : out <= 12'b000100100000;
501 : out <= 12'b000100011001;
502 : out <= 12'b000100011001;
503 : out <= 12'b000100011001;
504 : out <= 12'b000100011001;
505 : out <= 12'b000100011000;
506 : out <= 12'b000100011000;
507 : out <= 12'b000100011000;
508 : out <= 12'b000100011000;
509 : out <= 12'b000100010111;
510 : out <= 12'b000100010111;
511 : out <= 12'b000100010111;
512 : out <= 12'b000100010111;
513 : out <= 12'b000100010110;
514 : out <= 12'b000100010110;
515 : out <= 12'b000100010110;
516 : out <= 12'b000100010110;
517 : out <= 12'b000100010110;
518 : out <= 12'b000100010101;
519 : out <= 12'b000100010101;
520 : out <= 12'b000100010101;
521 : out <= 12'b000100010101;
522 : out <= 12'b000100010100;
523 : out <= 12'b000100010100;
524 : out <= 12'b000100010100;
525 : out <= 12'b000100010100;
526 : out <= 12'b000100010100;
527 : out <= 12'b000100010011;
528 : out <= 12'b000100010011;
529 : out <= 12'b000100010011;
530 : out <= 12'b000100010011;
531 : out <= 12'b000100010010;
532 : out <= 12'b000100010010;
533 : out <= 12'b000100010010;
534 : out <= 12'b000100010010;
535 : out <= 12'b000100010010;
536 : out <= 12'b000100010001;
537 : out <= 12'b000100010001;
538 : out <= 12'b000100010001;
539 : out <= 12'b000100010001;
540 : out <= 12'b000100010001;
541 : out <= 12'b000100010000;
542 : out <= 12'b000100010000;
543 : out <= 12'b000100010000;
544 : out <= 12'b000100010000;
545 : out <= 12'b000100010000;
546 : out <= 12'b000100001001;
547 : out <= 12'b000100001001;
548 : out <= 12'b000100001001;
549 : out <= 12'b000100001001;
550 : out <= 12'b000100001001;
551 : out <= 12'b000100001000;
552 : out <= 12'b000100001000;
553 : out <= 12'b000100001000;
554 : out <= 12'b000100001000;
555 : out <= 12'b000100001000;
556 : out <= 12'b000100000111;
557 : out <= 12'b000100000111;
558 : out <= 12'b000100000111;
559 : out <= 12'b000100000111;
560 : out <= 12'b000100000111;
561 : out <= 12'b000100000110;
562 : out <= 12'b000100000110;
563 : out <= 12'b000100000110;
564 : out <= 12'b000100000110;
565 : out <= 12'b000100000110;
566 : out <= 12'b000100000110;
567 : out <= 12'b000100000101;
568 : out <= 12'b000100000101;
569 : out <= 12'b000100000101;
570 : out <= 12'b000100000101;
571 : out <= 12'b000100000101;
572 : out <= 12'b000100000100;
573 : out <= 12'b000100000100;
574 : out <= 12'b000100000100;
575 : out <= 12'b000100000100;
576 : out <= 12'b000100000100;
577 : out <= 12'b000100000011;
578 : out <= 12'b000100000011;
579 : out <= 12'b000100000011;
580 : out <= 12'b000100000011;
581 : out <= 12'b000100000011;
582 : out <= 12'b000100000011;
583 : out <= 12'b000100000010;
584 : out <= 12'b000100000010;
585 : out <= 12'b000100000010;
586 : out <= 12'b000100000010;
587 : out <= 12'b000100000010;
588 : out <= 12'b000100000010;
589 : out <= 12'b000100000001;
590 : out <= 12'b000100000001;
591 : out <= 12'b000100000001;
592 : out <= 12'b000100000001;
593 : out <= 12'b000100000001;
594 : out <= 12'b000100000001;
595 : out <= 12'b000100000000;
596 : out <= 12'b000100000000;
597 : out <= 12'b000100000000;
598 : out <= 12'b000100000000;
599 : out <= 12'b000100000000;
600 : out <= 12'b000100000000;
601 : out <= 12'b000010011001;
602 : out <= 12'b000010011001;
603 : out <= 12'b000010011001;
604 : out <= 12'b000010011001;
605 : out <= 12'b000010011001;
606 : out <= 12'b000010011001;
607 : out <= 12'b000010011000;
608 : out <= 12'b000010011000;
609 : out <= 12'b000010011000;
610 : out <= 12'b000010011000;
611 : out <= 12'b000010011000;
612 : out <= 12'b000010011000;
613 : out <= 12'b000010010111;
614 : out <= 12'b000010010111;
615 : out <= 12'b000010010111;
616 : out <= 12'b000010010111;
617 : out <= 12'b000010010111;
618 : out <= 12'b000010010111;
619 : out <= 12'b000010010110;
620 : out <= 12'b000010010110;
621 : out <= 12'b000010010110;
622 : out <= 12'b000010010110;
623 : out <= 12'b000010010110;
624 : out <= 12'b000010010110;
625 : out <= 12'b000010010110;
626 : out <= 12'b000010010101;
627 : out <= 12'b000010010101;
628 : out <= 12'b000010010101;
629 : out <= 12'b000010010101;
630 : out <= 12'b000010010101;
631 : out <= 12'b000010010101;
632 : out <= 12'b000010010100;
633 : out <= 12'b000010010100;
634 : out <= 12'b000010010100;
635 : out <= 12'b000010010100;
636 : out <= 12'b000010010100;
637 : out <= 12'b000010010100;
638 : out <= 12'b000010010100;
639 : out <= 12'b000010010011;
640 : out <= 12'b000010010011;
641 : out <= 12'b000010010011;
642 : out <= 12'b000010010011;
643 : out <= 12'b000010010011;
644 : out <= 12'b000010010011;
645 : out <= 12'b000010010011;
646 : out <= 12'b000010010010;
647 : out <= 12'b000010010010;
648 : out <= 12'b000010010010;
649 : out <= 12'b000010010010;
650 : out <= 12'b000010010010;
651 : out <= 12'b000010010010;
652 : out <= 12'b000010010010;
653 : out <= 12'b000010010001;
654 : out <= 12'b000010010001;
655 : out <= 12'b000010010001;
656 : out <= 12'b000010010001;
657 : out <= 12'b000010010001;
658 : out <= 12'b000010010001;
659 : out <= 12'b000010010001;
660 : out <= 12'b000010010000;
661 : out <= 12'b000010010000;
662 : out <= 12'b000010010000;
663 : out <= 12'b000010010000;
664 : out <= 12'b000010010000;
665 : out <= 12'b000010010000;
666 : out <= 12'b000010010000;
667 : out <= 12'b000010001001;
668 : out <= 12'b000010001001;
669 : out <= 12'b000010001001;
670 : out <= 12'b000010001001;
671 : out <= 12'b000010001001;
672 : out <= 12'b000010001001;
673 : out <= 12'b000010001001;
674 : out <= 12'b000010001001;
675 : out <= 12'b000010001000;
676 : out <= 12'b000010001000;
677 : out <= 12'b000010001000;
678 : out <= 12'b000010001000;
679 : out <= 12'b000010001000;
680 : out <= 12'b000010001000;
681 : out <= 12'b000010001000;
682 : out <= 12'b000010000111;
683 : out <= 12'b000010000111;
684 : out <= 12'b000010000111;
685 : out <= 12'b000010000111;
686 : out <= 12'b000010000111;
687 : out <= 12'b000010000111;
688 : out <= 12'b000010000111;
689 : out <= 12'b000010000111;
690 : out <= 12'b000010000110;
691 : out <= 12'b000010000110;
692 : out <= 12'b000010000110;
693 : out <= 12'b000010000110;
694 : out <= 12'b000010000110;
695 : out <= 12'b000010000110;
696 : out <= 12'b000010000110;
697 : out <= 12'b000010000110;
698 : out <= 12'b000010000101;
699 : out <= 12'b000010000101;
700 : out <= 12'b000010000101;
701 : out <= 12'b000010000101;
702 : out <= 12'b000010000101;
703 : out <= 12'b000010000101;
704 : out <= 12'b000010000101;
705 : out <= 12'b000010000101;
706 : out <= 12'b000010000100;
707 : out <= 12'b000010000100;
708 : out <= 12'b000010000100;
709 : out <= 12'b000010000100;
710 : out <= 12'b000010000100;
711 : out <= 12'b000010000100;
712 : out <= 12'b000010000100;
713 : out <= 12'b000010000100;
714 : out <= 12'b000010000100;
715 : out <= 12'b000010000011;
716 : out <= 12'b000010000011;
717 : out <= 12'b000010000011;
718 : out <= 12'b000010000011;
719 : out <= 12'b000010000011;
720 : out <= 12'b000010000011;
721 : out <= 12'b000010000011;
722 : out <= 12'b000010000011;
723 : out <= 12'b000010000010;
724 : out <= 12'b000010000010;
725 : out <= 12'b000010000010;
726 : out <= 12'b000010000010;
727 : out <= 12'b000010000010;
728 : out <= 12'b000010000010;
729 : out <= 12'b000010000010;
730 : out <= 12'b000010000010;
731 : out <= 12'b000010000010;
732 : out <= 12'b000010000001;
733 : out <= 12'b000010000001;
734 : out <= 12'b000010000001;
735 : out <= 12'b000010000001;
736 : out <= 12'b000010000001;
737 : out <= 12'b000010000001;
738 : out <= 12'b000010000001;
739 : out <= 12'b000010000001;
740 : out <= 12'b000010000001;
741 : out <= 12'b000010000000;
742 : out <= 12'b000010000000;
743 : out <= 12'b000010000000;
744 : out <= 12'b000010000000;
745 : out <= 12'b000010000000;
746 : out <= 12'b000010000000;
747 : out <= 12'b000010000000;
748 : out <= 12'b000010000000;
749 : out <= 12'b000010000000;
750 : out <= 12'b000010000000;
751 : out <= 12'b000001111001;
752 : out <= 12'b000001111001;
753 : out <= 12'b000001111001;
754 : out <= 12'b000001111001;
755 : out <= 12'b000001111001;
756 : out <= 12'b000001111001;
757 : out <= 12'b000001111001;
758 : out <= 12'b000001111001;
759 : out <= 12'b000001111001;
760 : out <= 12'b000001111000;
761 : out <= 12'b000001111000;
762 : out <= 12'b000001111000;
763 : out <= 12'b000001111000;
764 : out <= 12'b000001111000;
765 : out <= 12'b000001111000;
766 : out <= 12'b000001111000;
767 : out <= 12'b000001111000;
768 : out <= 12'b000001111000;
769 : out <= 12'b000001111000;
770 : out <= 12'b000001110111;
771 : out <= 12'b000001110111;
772 : out <= 12'b000001110111;
773 : out <= 12'b000001110111;
774 : out <= 12'b000001110111;
775 : out <= 12'b000001110111;
776 : out <= 12'b000001110111;
777 : out <= 12'b000001110111;
778 : out <= 12'b000001110111;
779 : out <= 12'b000001110111;
780 : out <= 12'b000001110110;
781 : out <= 12'b000001110110;
782 : out <= 12'b000001110110;
783 : out <= 12'b000001110110;
784 : out <= 12'b000001110110;
785 : out <= 12'b000001110110;
786 : out <= 12'b000001110110;
787 : out <= 12'b000001110110;
788 : out <= 12'b000001110110;
789 : out <= 12'b000001110110;
790 : out <= 12'b000001110101;
791 : out <= 12'b000001110101;
792 : out <= 12'b000001110101;
793 : out <= 12'b000001110101;
794 : out <= 12'b000001110101;
795 : out <= 12'b000001110101;
796 : out <= 12'b000001110101;
797 : out <= 12'b000001110101;
798 : out <= 12'b000001110101;
799 : out <= 12'b000001110101;
800 : out <= 12'b000001110101;
801 : out <= 12'b000001110100;
802 : out <= 12'b000001110100;
803 : out <= 12'b000001110100;
804 : out <= 12'b000001110100;
805 : out <= 12'b000001110100;
806 : out <= 12'b000001110100;
807 : out <= 12'b000001110100;
808 : out <= 12'b000001110100;
809 : out <= 12'b000001110100;
810 : out <= 12'b000001110100;
811 : out <= 12'b000001110011;
812 : out <= 12'b000001110011;
813 : out <= 12'b000001110011;
814 : out <= 12'b000001110011;
815 : out <= 12'b000001110011;
816 : out <= 12'b000001110011;
817 : out <= 12'b000001110011;
818 : out <= 12'b000001110011;
819 : out <= 12'b000001110011;
820 : out <= 12'b000001110011;
821 : out <= 12'b000001110011;
822 : out <= 12'b000001110010;
823 : out <= 12'b000001110010;
824 : out <= 12'b000001110010;
825 : out <= 12'b000001110010;
826 : out <= 12'b000001110010;
827 : out <= 12'b000001110010;
828 : out <= 12'b000001110010;
829 : out <= 12'b000001110010;
830 : out <= 12'b000001110010;
831 : out <= 12'b000001110010;
832 : out <= 12'b000001110010;
833 : out <= 12'b000001110010;
834 : out <= 12'b000001110001;
835 : out <= 12'b000001110001;
836 : out <= 12'b000001110001;
837 : out <= 12'b000001110001;
838 : out <= 12'b000001110001;
839 : out <= 12'b000001110001;
840 : out <= 12'b000001110001;
841 : out <= 12'b000001110001;
842 : out <= 12'b000001110001;
843 : out <= 12'b000001110001;
844 : out <= 12'b000001110001;
845 : out <= 12'b000001110001;
846 : out <= 12'b000001110000;
847 : out <= 12'b000001110000;
848 : out <= 12'b000001110000;
849 : out <= 12'b000001110000;
850 : out <= 12'b000001110000;
851 : out <= 12'b000001110000;
852 : out <= 12'b000001110000;
853 : out <= 12'b000001110000;
854 : out <= 12'b000001110000;
855 : out <= 12'b000001110000;
856 : out <= 12'b000001110000;
857 : out <= 12'b000001110000;
858 : out <= 12'b000001101001;
859 : out <= 12'b000001101001;
860 : out <= 12'b000001101001;
861 : out <= 12'b000001101001;
862 : out <= 12'b000001101001;
863 : out <= 12'b000001101001;
864 : out <= 12'b000001101001;
865 : out <= 12'b000001101001;
866 : out <= 12'b000001101001;
867 : out <= 12'b000001101001;
868 : out <= 12'b000001101001;
869 : out <= 12'b000001101001;
870 : out <= 12'b000001101000;
871 : out <= 12'b000001101000;
872 : out <= 12'b000001101000;
873 : out <= 12'b000001101000;
874 : out <= 12'b000001101000;
875 : out <= 12'b000001101000;
876 : out <= 12'b000001101000;
877 : out <= 12'b000001101000;
878 : out <= 12'b000001101000;
879 : out <= 12'b000001101000;
880 : out <= 12'b000001101000;
881 : out <= 12'b000001101000;
882 : out <= 12'b000001101000;
883 : out <= 12'b000001100111;
884 : out <= 12'b000001100111;
885 : out <= 12'b000001100111;
886 : out <= 12'b000001100111;
887 : out <= 12'b000001100111;
888 : out <= 12'b000001100111;
889 : out <= 12'b000001100111;
890 : out <= 12'b000001100111;
891 : out <= 12'b000001100111;
892 : out <= 12'b000001100111;
893 : out <= 12'b000001100111;
894 : out <= 12'b000001100111;
895 : out <= 12'b000001100111;
896 : out <= 12'b000001100110;
897 : out <= 12'b000001100110;
898 : out <= 12'b000001100110;
899 : out <= 12'b000001100110;
900 : out <= 12'b000001100110;
901 : out <= 12'b000001100110;
902 : out <= 12'b000001100110;
903 : out <= 12'b000001100110;
904 : out <= 12'b000001100110;
905 : out <= 12'b000001100110;
906 : out <= 12'b000001100110;
907 : out <= 12'b000001100110;
908 : out <= 12'b000001100110;
909 : out <= 12'b000001100110;
910 : out <= 12'b000001100101;
911 : out <= 12'b000001100101;
912 : out <= 12'b000001100101;
913 : out <= 12'b000001100101;
914 : out <= 12'b000001100101;
915 : out <= 12'b000001100101;
916 : out <= 12'b000001100101;
917 : out <= 12'b000001100101;
918 : out <= 12'b000001100101;
919 : out <= 12'b000001100101;
920 : out <= 12'b000001100101;
921 : out <= 12'b000001100101;
922 : out <= 12'b000001100101;
923 : out <= 12'b000001100101;
924 : out <= 12'b000001100100;
925 : out <= 12'b000001100100;
926 : out <= 12'b000001100100;
927 : out <= 12'b000001100100;
928 : out <= 12'b000001100100;
929 : out <= 12'b000001100100;
930 : out <= 12'b000001100100;
931 : out <= 12'b000001100100;
932 : out <= 12'b000001100100;
933 : out <= 12'b000001100100;
934 : out <= 12'b000001100100;
935 : out <= 12'b000001100100;
936 : out <= 12'b000001100100;
937 : out <= 12'b000001100100;
938 : out <= 12'b000001100011;
939 : out <= 12'b000001100011;
940 : out <= 12'b000001100011;
941 : out <= 12'b000001100011;
942 : out <= 12'b000001100011;
943 : out <= 12'b000001100011;
944 : out <= 12'b000001100011;
945 : out <= 12'b000001100011;
946 : out <= 12'b000001100011;
947 : out <= 12'b000001100011;
948 : out <= 12'b000001100011;
949 : out <= 12'b000001100011;
950 : out <= 12'b000001100011;
951 : out <= 12'b000001100011;
952 : out <= 12'b000001100011;
953 : out <= 12'b000001100010;
954 : out <= 12'b000001100010;
955 : out <= 12'b000001100010;
956 : out <= 12'b000001100010;
957 : out <= 12'b000001100010;
958 : out <= 12'b000001100010;
959 : out <= 12'b000001100010;
960 : out <= 12'b000001100010;
961 : out <= 12'b000001100010;
962 : out <= 12'b000001100010;
963 : out <= 12'b000001100010;
964 : out <= 12'b000001100010;
965 : out <= 12'b000001100010;
966 : out <= 12'b000001100010;
967 : out <= 12'b000001100010;
968 : out <= 12'b000001100001;
969 : out <= 12'b000001100001;
970 : out <= 12'b000001100001;
971 : out <= 12'b000001100001;
972 : out <= 12'b000001100001;
973 : out <= 12'b000001100001;
974 : out <= 12'b000001100001;
975 : out <= 12'b000001100001;
976 : out <= 12'b000001100001;
977 : out <= 12'b000001100001;
978 : out <= 12'b000001100001;
979 : out <= 12'b000001100001;
980 : out <= 12'b000001100001;
981 : out <= 12'b000001100001;
982 : out <= 12'b000001100001;
983 : out <= 12'b000001100001;
984 : out <= 12'b000001100000;
985 : out <= 12'b000001100000;
986 : out <= 12'b000001100000;
987 : out <= 12'b000001100000;
988 : out <= 12'b000001100000;
989 : out <= 12'b000001100000;
990 : out <= 12'b000001100000;
991 : out <= 12'b000001100000;
992 : out <= 12'b000001100000;
993 : out <= 12'b000001100000;
994 : out <= 12'b000001100000;
995 : out <= 12'b000001100000;
996 : out <= 12'b000001100000;
997 : out <= 12'b000001100000;
998 : out <= 12'b000001100000;
999 : out <= 12'b000001100000;
1000 : out <= 12'b000001100000;
1001 : out <= 12'b000001011001;
1002 : out <= 12'b000001011001;
1003 : out <= 12'b000001011001;
1004 : out <= 12'b000001011001;
1005 : out <= 12'b000001011001;
1006 : out <= 12'b000001011001;
1007 : out <= 12'b000001011001;
1008 : out <= 12'b000001011001;
1009 : out <= 12'b000001011001;
1010 : out <= 12'b000001011001;
1011 : out <= 12'b000001011001;
1012 : out <= 12'b000001011001;
1013 : out <= 12'b000001011001;
1014 : out <= 12'b000001011001;
1015 : out <= 12'b000001011001;
1016 : out <= 12'b000001011001;
1017 : out <= 12'b000001011000;
1018 : out <= 12'b000001011000;
1019 : out <= 12'b000001011000;
1020 : out <= 12'b000001011000;
1021 : out <= 12'b000001011000;
1022 : out <= 12'b000001011000;
1023 : out <= 12'b000001011000;
1024 : out <= 12'b000001011000;
1025 : out <= 12'b000001011000;
1026 : out <= 12'b000001011000;
1027 : out <= 12'b000001011000;
1028 : out <= 12'b000001011000;
1029 : out <= 12'b000001011000;
1030 : out <= 12'b000001011000;
1031 : out <= 12'b000001011000;
1032 : out <= 12'b000001011000;
1033 : out <= 12'b000001011000;
1034 : out <= 12'b000001011000;
1035 : out <= 12'b000001010111;
1036 : out <= 12'b000001010111;
1037 : out <= 12'b000001010111;
1038 : out <= 12'b000001010111;
1039 : out <= 12'b000001010111;
1040 : out <= 12'b000001010111;
1041 : out <= 12'b000001010111;
1042 : out <= 12'b000001010111;
1043 : out <= 12'b000001010111;
1044 : out <= 12'b000001010111;
1045 : out <= 12'b000001010111;
1046 : out <= 12'b000001010111;
1047 : out <= 12'b000001010111;
1048 : out <= 12'b000001010111;
1049 : out <= 12'b000001010111;
1050 : out <= 12'b000001010111;
1051 : out <= 12'b000001010111;
1052 : out <= 12'b000001010111;
1053 : out <= 12'b000001010110;
1054 : out <= 12'b000001010110;
1055 : out <= 12'b000001010110;
1056 : out <= 12'b000001010110;
1057 : out <= 12'b000001010110;
1058 : out <= 12'b000001010110;
1059 : out <= 12'b000001010110;
1060 : out <= 12'b000001010110;
1061 : out <= 12'b000001010110;
1062 : out <= 12'b000001010110;
1063 : out <= 12'b000001010110;
1064 : out <= 12'b000001010110;
1065 : out <= 12'b000001010110;
1066 : out <= 12'b000001010110;
1067 : out <= 12'b000001010110;
1068 : out <= 12'b000001010110;
1069 : out <= 12'b000001010110;
1070 : out <= 12'b000001010110;
1071 : out <= 12'b000001010110;
1072 : out <= 12'b000001010101;
1073 : out <= 12'b000001010101;
1074 : out <= 12'b000001010101;
1075 : out <= 12'b000001010101;
1076 : out <= 12'b000001010101;
1077 : out <= 12'b000001010101;
1078 : out <= 12'b000001010101;
1079 : out <= 12'b000001010101;
1080 : out <= 12'b000001010101;
1081 : out <= 12'b000001010101;
1082 : out <= 12'b000001010101;
1083 : out <= 12'b000001010101;
1084 : out <= 12'b000001010101;
1085 : out <= 12'b000001010101;
1086 : out <= 12'b000001010101;
1087 : out <= 12'b000001010101;
1088 : out <= 12'b000001010101;
1089 : out <= 12'b000001010101;
1090 : out <= 12'b000001010101;
1091 : out <= 12'b000001010100;
1092 : out <= 12'b000001010100;
1093 : out <= 12'b000001010100;
1094 : out <= 12'b000001010100;
1095 : out <= 12'b000001010100;
1096 : out <= 12'b000001010100;
1097 : out <= 12'b000001010100;
1098 : out <= 12'b000001010100;
1099 : out <= 12'b000001010100;
1100 : out <= 12'b000001010100;
1101 : out <= 12'b000001010100;
1102 : out <= 12'b000001010100;
1103 : out <= 12'b000001010100;
1104 : out <= 12'b000001010100;
1105 : out <= 12'b000001010100;
1106 : out <= 12'b000001010100;
1107 : out <= 12'b000001010100;
1108 : out <= 12'b000001010100;
1109 : out <= 12'b000001010100;
1110 : out <= 12'b000001010100;
1111 : out <= 12'b000001010100;
1112 : out <= 12'b000001010011;
1113 : out <= 12'b000001010011;
1114 : out <= 12'b000001010011;
1115 : out <= 12'b000001010011;
1116 : out <= 12'b000001010011;
1117 : out <= 12'b000001010011;
1118 : out <= 12'b000001010011;
1119 : out <= 12'b000001010011;
1120 : out <= 12'b000001010011;
1121 : out <= 12'b000001010011;
1122 : out <= 12'b000001010011;
1123 : out <= 12'b000001010011;
1124 : out <= 12'b000001010011;
1125 : out <= 12'b000001010011;
1126 : out <= 12'b000001010011;
1127 : out <= 12'b000001010011;
1128 : out <= 12'b000001010011;
1129 : out <= 12'b000001010011;
1130 : out <= 12'b000001010011;
1131 : out <= 12'b000001010011;
1132 : out <= 12'b000001010011;
1133 : out <= 12'b000001010010;
1134 : out <= 12'b000001010010;
1135 : out <= 12'b000001010010;
1136 : out <= 12'b000001010010;
1137 : out <= 12'b000001010010;
1138 : out <= 12'b000001010010;
1139 : out <= 12'b000001010010;
1140 : out <= 12'b000001010010;
1141 : out <= 12'b000001010010;
1142 : out <= 12'b000001010010;
1143 : out <= 12'b000001010010;
1144 : out <= 12'b000001010010;
1145 : out <= 12'b000001010010;
1146 : out <= 12'b000001010010;
1147 : out <= 12'b000001010010;
1148 : out <= 12'b000001010010;
1149 : out <= 12'b000001010010;
1150 : out <= 12'b000001010010;
1151 : out <= 12'b000001010010;
1152 : out <= 12'b000001010010;
1153 : out <= 12'b000001010010;
1154 : out <= 12'b000001010001;
1155 : out <= 12'b000001010001;
1156 : out <= 12'b000001010001;
1157 : out <= 12'b000001010001;
1158 : out <= 12'b000001010001;
1159 : out <= 12'b000001010001;
1160 : out <= 12'b000001010001;
1161 : out <= 12'b000001010001;
1162 : out <= 12'b000001010001;
1163 : out <= 12'b000001010001;
1164 : out <= 12'b000001010001;
1165 : out <= 12'b000001010001;
1166 : out <= 12'b000001010001;
1167 : out <= 12'b000001010001;
1168 : out <= 12'b000001010001;
1169 : out <= 12'b000001010001;
1170 : out <= 12'b000001010001;
1171 : out <= 12'b000001010001;
1172 : out <= 12'b000001010001;
1173 : out <= 12'b000001010001;
1174 : out <= 12'b000001010001;
1175 : out <= 12'b000001010001;
1176 : out <= 12'b000001010001;
1177 : out <= 12'b000001010000;
1178 : out <= 12'b000001010000;
1179 : out <= 12'b000001010000;
1180 : out <= 12'b000001010000;
1181 : out <= 12'b000001010000;
1182 : out <= 12'b000001010000;
1183 : out <= 12'b000001010000;
1184 : out <= 12'b000001010000;
1185 : out <= 12'b000001010000;
1186 : out <= 12'b000001010000;
1187 : out <= 12'b000001010000;
1188 : out <= 12'b000001010000;
1189 : out <= 12'b000001010000;
1190 : out <= 12'b000001010000;
1191 : out <= 12'b000001010000;
1192 : out <= 12'b000001010000;
1193 : out <= 12'b000001010000;
1194 : out <= 12'b000001010000;
1195 : out <= 12'b000001010000;
1196 : out <= 12'b000001010000;
1197 : out <= 12'b000001010000;
1198 : out <= 12'b000001010000;
1199 : out <= 12'b000001010000;
1200 : out <= 12'b000001010000;
1201 : out <= 12'b000001001001;
1202 : out <= 12'b000001001001;
1203 : out <= 12'b000001001001;
1204 : out <= 12'b000001001001;
1205 : out <= 12'b000001001001;
1206 : out <= 12'b000001001001;
1207 : out <= 12'b000001001001;
1208 : out <= 12'b000001001001;
1209 : out <= 12'b000001001001;
1210 : out <= 12'b000001001001;
1211 : out <= 12'b000001001001;
1212 : out <= 12'b000001001001;
1213 : out <= 12'b000001001001;
1214 : out <= 12'b000001001001;
1215 : out <= 12'b000001001001;
1216 : out <= 12'b000001001001;
1217 : out <= 12'b000001001001;
1218 : out <= 12'b000001001001;
1219 : out <= 12'b000001001001;
1220 : out <= 12'b000001001001;
1221 : out <= 12'b000001001001;
1222 : out <= 12'b000001001001;
1223 : out <= 12'b000001001001;
1224 : out <= 12'b000001001001;
1225 : out <= 12'b000001001000;
1226 : out <= 12'b000001001000;
1227 : out <= 12'b000001001000;
1228 : out <= 12'b000001001000;
1229 : out <= 12'b000001001000;
1230 : out <= 12'b000001001000;
1231 : out <= 12'b000001001000;
1232 : out <= 12'b000001001000;
1233 : out <= 12'b000001001000;
1234 : out <= 12'b000001001000;
1235 : out <= 12'b000001001000;
1236 : out <= 12'b000001001000;
1237 : out <= 12'b000001001000;
1238 : out <= 12'b000001001000;
1239 : out <= 12'b000001001000;
1240 : out <= 12'b000001001000;
1241 : out <= 12'b000001001000;
1242 : out <= 12'b000001001000;
1243 : out <= 12'b000001001000;
1244 : out <= 12'b000001001000;
1245 : out <= 12'b000001001000;
1246 : out <= 12'b000001001000;
1247 : out <= 12'b000001001000;
1248 : out <= 12'b000001001000;
1249 : out <= 12'b000001001000;
1250 : out <= 12'b000001001000;
1251 : out <= 12'b000001000111;
1252 : out <= 12'b000001000111;
1253 : out <= 12'b000001000111;
1254 : out <= 12'b000001000111;
1255 : out <= 12'b000001000111;
1256 : out <= 12'b000001000111;
1257 : out <= 12'b000001000111;
1258 : out <= 12'b000001000111;
1259 : out <= 12'b000001000111;
1260 : out <= 12'b000001000111;
1261 : out <= 12'b000001000111;
1262 : out <= 12'b000001000111;
1263 : out <= 12'b000001000111;
1264 : out <= 12'b000001000111;
1265 : out <= 12'b000001000111;
1266 : out <= 12'b000001000111;
1267 : out <= 12'b000001000111;
1268 : out <= 12'b000001000111;
1269 : out <= 12'b000001000111;
1270 : out <= 12'b000001000111;
1271 : out <= 12'b000001000111;
1272 : out <= 12'b000001000111;
1273 : out <= 12'b000001000111;
1274 : out <= 12'b000001000111;
1275 : out <= 12'b000001000111;
1276 : out <= 12'b000001000111;
1277 : out <= 12'b000001000110;
1278 : out <= 12'b000001000110;
1279 : out <= 12'b000001000110;
1280 : out <= 12'b000001000110;
1281 : out <= 12'b000001000110;
1282 : out <= 12'b000001000110;
1283 : out <= 12'b000001000110;
1284 : out <= 12'b000001000110;
1285 : out <= 12'b000001000110;
1286 : out <= 12'b000001000110;
1287 : out <= 12'b000001000110;
1288 : out <= 12'b000001000110;
1289 : out <= 12'b000001000110;
1290 : out <= 12'b000001000110;
1291 : out <= 12'b000001000110;
1292 : out <= 12'b000001000110;
1293 : out <= 12'b000001000110;
1294 : out <= 12'b000001000110;
1295 : out <= 12'b000001000110;
1296 : out <= 12'b000001000110;
1297 : out <= 12'b000001000110;
1298 : out <= 12'b000001000110;
1299 : out <= 12'b000001000110;
1300 : out <= 12'b000001000110;
1301 : out <= 12'b000001000110;
1302 : out <= 12'b000001000110;
1303 : out <= 12'b000001000110;
1304 : out <= 12'b000001000110;
1305 : out <= 12'b000001000101;
1306 : out <= 12'b000001000101;
1307 : out <= 12'b000001000101;
1308 : out <= 12'b000001000101;
1309 : out <= 12'b000001000101;
1310 : out <= 12'b000001000101;
1311 : out <= 12'b000001000101;
1312 : out <= 12'b000001000101;
1313 : out <= 12'b000001000101;
1314 : out <= 12'b000001000101;
1315 : out <= 12'b000001000101;
1316 : out <= 12'b000001000101;
1317 : out <= 12'b000001000101;
1318 : out <= 12'b000001000101;
1319 : out <= 12'b000001000101;
1320 : out <= 12'b000001000101;
1321 : out <= 12'b000001000101;
1322 : out <= 12'b000001000101;
1323 : out <= 12'b000001000101;
1324 : out <= 12'b000001000101;
1325 : out <= 12'b000001000101;
1326 : out <= 12'b000001000101;
1327 : out <= 12'b000001000101;
1328 : out <= 12'b000001000101;
1329 : out <= 12'b000001000101;
1330 : out <= 12'b000001000101;
1331 : out <= 12'b000001000101;
1332 : out <= 12'b000001000101;
1333 : out <= 12'b000001000101;
1334 : out <= 12'b000001000100;
1335 : out <= 12'b000001000100;
1336 : out <= 12'b000001000100;
1337 : out <= 12'b000001000100;
1338 : out <= 12'b000001000100;
1339 : out <= 12'b000001000100;
1340 : out <= 12'b000001000100;
1341 : out <= 12'b000001000100;
1342 : out <= 12'b000001000100;
1343 : out <= 12'b000001000100;
1344 : out <= 12'b000001000100;
1345 : out <= 12'b000001000100;
1346 : out <= 12'b000001000100;
1347 : out <= 12'b000001000100;
1348 : out <= 12'b000001000100;
1349 : out <= 12'b000001000100;
1350 : out <= 12'b000001000100;
1351 : out <= 12'b000001000100;
1352 : out <= 12'b000001000100;
1353 : out <= 12'b000001000100;
1354 : out <= 12'b000001000100;
1355 : out <= 12'b000001000100;
1356 : out <= 12'b000001000100;
1357 : out <= 12'b000001000100;
1358 : out <= 12'b000001000100;
1359 : out <= 12'b000001000100;
1360 : out <= 12'b000001000100;
1361 : out <= 12'b000001000100;
1362 : out <= 12'b000001000100;
1363 : out <= 12'b000001000100;
1364 : out <= 12'b000001000011;
1365 : out <= 12'b000001000011;
1366 : out <= 12'b000001000011;
1367 : out <= 12'b000001000011;
1368 : out <= 12'b000001000011;
1369 : out <= 12'b000001000011;
1370 : out <= 12'b000001000011;
1371 : out <= 12'b000001000011;
1372 : out <= 12'b000001000011;
1373 : out <= 12'b000001000011;
1374 : out <= 12'b000001000011;
1375 : out <= 12'b000001000011;
1376 : out <= 12'b000001000011;
1377 : out <= 12'b000001000011;
1378 : out <= 12'b000001000011;
1379 : out <= 12'b000001000011;
1380 : out <= 12'b000001000011;
1381 : out <= 12'b000001000011;
1382 : out <= 12'b000001000011;
1383 : out <= 12'b000001000011;
1384 : out <= 12'b000001000011;
1385 : out <= 12'b000001000011;
1386 : out <= 12'b000001000011;
1387 : out <= 12'b000001000011;
1388 : out <= 12'b000001000011;
1389 : out <= 12'b000001000011;
1390 : out <= 12'b000001000011;
1391 : out <= 12'b000001000011;
1392 : out <= 12'b000001000011;
1393 : out <= 12'b000001000011;
1394 : out <= 12'b000001000011;
1395 : out <= 12'b000001000011;
1396 : out <= 12'b000001000010;
1397 : out <= 12'b000001000010;
1398 : out <= 12'b000001000010;
1399 : out <= 12'b000001000010;
1400 : out <= 12'b000001000010;
1401 : out <= 12'b000001000010;
1402 : out <= 12'b000001000010;
1403 : out <= 12'b000001000010;
1404 : out <= 12'b000001000010;
1405 : out <= 12'b000001000010;
1406 : out <= 12'b000001000010;
1407 : out <= 12'b000001000010;
1408 : out <= 12'b000001000010;
1409 : out <= 12'b000001000010;
1410 : out <= 12'b000001000010;
1411 : out <= 12'b000001000010;
1412 : out <= 12'b000001000010;
1413 : out <= 12'b000001000010;
1414 : out <= 12'b000001000010;
1415 : out <= 12'b000001000010;
1416 : out <= 12'b000001000010;
1417 : out <= 12'b000001000010;
1418 : out <= 12'b000001000010;
1419 : out <= 12'b000001000010;
1420 : out <= 12'b000001000010;
1421 : out <= 12'b000001000010;
1422 : out <= 12'b000001000010;
1423 : out <= 12'b000001000010;
1424 : out <= 12'b000001000010;
1425 : out <= 12'b000001000010;
1426 : out <= 12'b000001000010;
1427 : out <= 12'b000001000010;
1428 : out <= 12'b000001000010;
1429 : out <= 12'b000001000001;
1430 : out <= 12'b000001000001;
1431 : out <= 12'b000001000001;
1432 : out <= 12'b000001000001;
1433 : out <= 12'b000001000001;
1434 : out <= 12'b000001000001;
1435 : out <= 12'b000001000001;
1436 : out <= 12'b000001000001;
1437 : out <= 12'b000001000001;
1438 : out <= 12'b000001000001;
1439 : out <= 12'b000001000001;
1440 : out <= 12'b000001000001;
1441 : out <= 12'b000001000001;
1442 : out <= 12'b000001000001;
1443 : out <= 12'b000001000001;
1444 : out <= 12'b000001000001;
1445 : out <= 12'b000001000001;
1446 : out <= 12'b000001000001;
1447 : out <= 12'b000001000001;
1448 : out <= 12'b000001000001;
1449 : out <= 12'b000001000001;
1450 : out <= 12'b000001000001;
1451 : out <= 12'b000001000001;
1452 : out <= 12'b000001000001;
1453 : out <= 12'b000001000001;
1454 : out <= 12'b000001000001;
1455 : out <= 12'b000001000001;
1456 : out <= 12'b000001000001;
1457 : out <= 12'b000001000001;
1458 : out <= 12'b000001000001;
1459 : out <= 12'b000001000001;
1460 : out <= 12'b000001000001;
1461 : out <= 12'b000001000001;
1462 : out <= 12'b000001000001;
1463 : out <= 12'b000001000001;
1464 : out <= 12'b000001000000;
1465 : out <= 12'b000001000000;
1466 : out <= 12'b000001000000;
1467 : out <= 12'b000001000000;
1468 : out <= 12'b000001000000;
1469 : out <= 12'b000001000000;
1470 : out <= 12'b000001000000;
1471 : out <= 12'b000001000000;
1472 : out <= 12'b000001000000;
1473 : out <= 12'b000001000000;
1474 : out <= 12'b000001000000;
1475 : out <= 12'b000001000000;
1476 : out <= 12'b000001000000;
1477 : out <= 12'b000001000000;
1478 : out <= 12'b000001000000;
1479 : out <= 12'b000001000000;
1480 : out <= 12'b000001000000;
1481 : out <= 12'b000001000000;
1482 : out <= 12'b000001000000;
1483 : out <= 12'b000001000000;
1484 : out <= 12'b000001000000;
1485 : out <= 12'b000001000000;
1486 : out <= 12'b000001000000;
1487 : out <= 12'b000001000000;
1488 : out <= 12'b000001000000;
1489 : out <= 12'b000001000000;
1490 : out <= 12'b000001000000;
1491 : out <= 12'b000001000000;
1492 : out <= 12'b000001000000;
1493 : out <= 12'b000001000000;
1494 : out <= 12'b000001000000;
1495 : out <= 12'b000001000000;
1496 : out <= 12'b000001000000;
1497 : out <= 12'b000001000000;
1498 : out <= 12'b000001000000;
1499 : out <= 12'b000001000000;
1500 : out <= 12'b000001000000;
1501 : out <= 12'b000000111001;
1502 : out <= 12'b000000111001;
1503 : out <= 12'b000000111001;
1504 : out <= 12'b000000111001;
1505 : out <= 12'b000000111001;
1506 : out <= 12'b000000111001;
1507 : out <= 12'b000000111001;
1508 : out <= 12'b000000111001;
1509 : out <= 12'b000000111001;
1510 : out <= 12'b000000111001;
1511 : out <= 12'b000000111001;
1512 : out <= 12'b000000111001;
1513 : out <= 12'b000000111001;
1514 : out <= 12'b000000111001;
1515 : out <= 12'b000000111001;
1516 : out <= 12'b000000111001;
1517 : out <= 12'b000000111001;
1518 : out <= 12'b000000111001;
1519 : out <= 12'b000000111001;
1520 : out <= 12'b000000111001;
1521 : out <= 12'b000000111001;
1522 : out <= 12'b000000111001;
1523 : out <= 12'b000000111001;
1524 : out <= 12'b000000111001;
1525 : out <= 12'b000000111001;
1526 : out <= 12'b000000111001;
1527 : out <= 12'b000000111001;
1528 : out <= 12'b000000111001;
1529 : out <= 12'b000000111001;
1530 : out <= 12'b000000111001;
1531 : out <= 12'b000000111001;
1532 : out <= 12'b000000111001;
1533 : out <= 12'b000000111001;
1534 : out <= 12'b000000111001;
1535 : out <= 12'b000000111001;
1536 : out <= 12'b000000111001;
1537 : out <= 12'b000000111001;
1538 : out <= 12'b000000111001;
1539 : out <= 12'b000000111000;
1540 : out <= 12'b000000111000;
1541 : out <= 12'b000000111000;
1542 : out <= 12'b000000111000;
1543 : out <= 12'b000000111000;
1544 : out <= 12'b000000111000;
1545 : out <= 12'b000000111000;
1546 : out <= 12'b000000111000;
1547 : out <= 12'b000000111000;
1548 : out <= 12'b000000111000;
1549 : out <= 12'b000000111000;
1550 : out <= 12'b000000111000;
1551 : out <= 12'b000000111000;
1552 : out <= 12'b000000111000;
1553 : out <= 12'b000000111000;
1554 : out <= 12'b000000111000;
1555 : out <= 12'b000000111000;
1556 : out <= 12'b000000111000;
1557 : out <= 12'b000000111000;
1558 : out <= 12'b000000111000;
1559 : out <= 12'b000000111000;
1560 : out <= 12'b000000111000;
1561 : out <= 12'b000000111000;
1562 : out <= 12'b000000111000;
1563 : out <= 12'b000000111000;
1564 : out <= 12'b000000111000;
1565 : out <= 12'b000000111000;
1566 : out <= 12'b000000111000;
1567 : out <= 12'b000000111000;
1568 : out <= 12'b000000111000;
1569 : out <= 12'b000000111000;
1570 : out <= 12'b000000111000;
1571 : out <= 12'b000000111000;
1572 : out <= 12'b000000111000;
1573 : out <= 12'b000000111000;
1574 : out <= 12'b000000111000;
1575 : out <= 12'b000000111000;
1576 : out <= 12'b000000111000;
1577 : out <= 12'b000000111000;
1578 : out <= 12'b000000111000;
1579 : out <= 12'b000000110111;
1580 : out <= 12'b000000110111;
1581 : out <= 12'b000000110111;
1582 : out <= 12'b000000110111;
1583 : out <= 12'b000000110111;
1584 : out <= 12'b000000110111;
1585 : out <= 12'b000000110111;
1586 : out <= 12'b000000110111;
1587 : out <= 12'b000000110111;
1588 : out <= 12'b000000110111;
1589 : out <= 12'b000000110111;
1590 : out <= 12'b000000110111;
1591 : out <= 12'b000000110111;
1592 : out <= 12'b000000110111;
1593 : out <= 12'b000000110111;
1594 : out <= 12'b000000110111;
1595 : out <= 12'b000000110111;
1596 : out <= 12'b000000110111;
1597 : out <= 12'b000000110111;
1598 : out <= 12'b000000110111;
1599 : out <= 12'b000000110111;
1600 : out <= 12'b000000110111;
1601 : out <= 12'b000000110111;
1602 : out <= 12'b000000110111;
1603 : out <= 12'b000000110111;
1604 : out <= 12'b000000110111;
1605 : out <= 12'b000000110111;
1606 : out <= 12'b000000110111;
1607 : out <= 12'b000000110111;
1608 : out <= 12'b000000110111;
1609 : out <= 12'b000000110111;
1610 : out <= 12'b000000110111;
1611 : out <= 12'b000000110111;
1612 : out <= 12'b000000110111;
1613 : out <= 12'b000000110111;
1614 : out <= 12'b000000110111;
1615 : out <= 12'b000000110111;
1616 : out <= 12'b000000110111;
1617 : out <= 12'b000000110111;
1618 : out <= 12'b000000110111;
1619 : out <= 12'b000000110111;
1620 : out <= 12'b000000110111;
1621 : out <= 12'b000000110111;
1622 : out <= 12'b000000110110;
1623 : out <= 12'b000000110110;
1624 : out <= 12'b000000110110;
1625 : out <= 12'b000000110110;
1626 : out <= 12'b000000110110;
1627 : out <= 12'b000000110110;
1628 : out <= 12'b000000110110;
1629 : out <= 12'b000000110110;
1630 : out <= 12'b000000110110;
1631 : out <= 12'b000000110110;
1632 : out <= 12'b000000110110;
1633 : out <= 12'b000000110110;
1634 : out <= 12'b000000110110;
1635 : out <= 12'b000000110110;
1636 : out <= 12'b000000110110;
1637 : out <= 12'b000000110110;
1638 : out <= 12'b000000110110;
1639 : out <= 12'b000000110110;
1640 : out <= 12'b000000110110;
1641 : out <= 12'b000000110110;
1642 : out <= 12'b000000110110;
1643 : out <= 12'b000000110110;
1644 : out <= 12'b000000110110;
1645 : out <= 12'b000000110110;
1646 : out <= 12'b000000110110;
1647 : out <= 12'b000000110110;
1648 : out <= 12'b000000110110;
1649 : out <= 12'b000000110110;
1650 : out <= 12'b000000110110;
1651 : out <= 12'b000000110110;
1652 : out <= 12'b000000110110;
1653 : out <= 12'b000000110110;
1654 : out <= 12'b000000110110;
1655 : out <= 12'b000000110110;
1656 : out <= 12'b000000110110;
1657 : out <= 12'b000000110110;
1658 : out <= 12'b000000110110;
1659 : out <= 12'b000000110110;
1660 : out <= 12'b000000110110;
1661 : out <= 12'b000000110110;
1662 : out <= 12'b000000110110;
1663 : out <= 12'b000000110110;
1664 : out <= 12'b000000110110;
1665 : out <= 12'b000000110110;
1666 : out <= 12'b000000110110;
1667 : out <= 12'b000000110101;
1668 : out <= 12'b000000110101;
1669 : out <= 12'b000000110101;
1670 : out <= 12'b000000110101;
1671 : out <= 12'b000000110101;
1672 : out <= 12'b000000110101;
1673 : out <= 12'b000000110101;
1674 : out <= 12'b000000110101;
1675 : out <= 12'b000000110101;
1676 : out <= 12'b000000110101;
1677 : out <= 12'b000000110101;
1678 : out <= 12'b000000110101;
1679 : out <= 12'b000000110101;
1680 : out <= 12'b000000110101;
1681 : out <= 12'b000000110101;
1682 : out <= 12'b000000110101;
1683 : out <= 12'b000000110101;
1684 : out <= 12'b000000110101;
1685 : out <= 12'b000000110101;
1686 : out <= 12'b000000110101;
1687 : out <= 12'b000000110101;
1688 : out <= 12'b000000110101;
1689 : out <= 12'b000000110101;
1690 : out <= 12'b000000110101;
1691 : out <= 12'b000000110101;
1692 : out <= 12'b000000110101;
1693 : out <= 12'b000000110101;
1694 : out <= 12'b000000110101;
1695 : out <= 12'b000000110101;
1696 : out <= 12'b000000110101;
1697 : out <= 12'b000000110101;
1698 : out <= 12'b000000110101;
1699 : out <= 12'b000000110101;
1700 : out <= 12'b000000110101;
1701 : out <= 12'b000000110101;
1702 : out <= 12'b000000110101;
1703 : out <= 12'b000000110101;
1704 : out <= 12'b000000110101;
1705 : out <= 12'b000000110101;
1706 : out <= 12'b000000110101;
1707 : out <= 12'b000000110101;
1708 : out <= 12'b000000110101;
1709 : out <= 12'b000000110101;
1710 : out <= 12'b000000110101;
1711 : out <= 12'b000000110101;
1712 : out <= 12'b000000110101;
1713 : out <= 12'b000000110101;
1714 : out <= 12'b000000110101;
1715 : out <= 12'b000000110100;
1716 : out <= 12'b000000110100;
1717 : out <= 12'b000000110100;
1718 : out <= 12'b000000110100;
1719 : out <= 12'b000000110100;
1720 : out <= 12'b000000110100;
1721 : out <= 12'b000000110100;
1722 : out <= 12'b000000110100;
1723 : out <= 12'b000000110100;
1724 : out <= 12'b000000110100;
1725 : out <= 12'b000000110100;
1726 : out <= 12'b000000110100;
1727 : out <= 12'b000000110100;
1728 : out <= 12'b000000110100;
1729 : out <= 12'b000000110100;
1730 : out <= 12'b000000110100;
1731 : out <= 12'b000000110100;
1732 : out <= 12'b000000110100;
1733 : out <= 12'b000000110100;
1734 : out <= 12'b000000110100;
1735 : out <= 12'b000000110100;
1736 : out <= 12'b000000110100;
1737 : out <= 12'b000000110100;
1738 : out <= 12'b000000110100;
1739 : out <= 12'b000000110100;
1740 : out <= 12'b000000110100;
1741 : out <= 12'b000000110100;
1742 : out <= 12'b000000110100;
1743 : out <= 12'b000000110100;
1744 : out <= 12'b000000110100;
1745 : out <= 12'b000000110100;
1746 : out <= 12'b000000110100;
1747 : out <= 12'b000000110100;
1748 : out <= 12'b000000110100;
1749 : out <= 12'b000000110100;
1750 : out <= 12'b000000110100;
1751 : out <= 12'b000000110100;
1752 : out <= 12'b000000110100;
1753 : out <= 12'b000000110100;
1754 : out <= 12'b000000110100;
1755 : out <= 12'b000000110100;
1756 : out <= 12'b000000110100;
1757 : out <= 12'b000000110100;
1758 : out <= 12'b000000110100;
1759 : out <= 12'b000000110100;
1760 : out <= 12'b000000110100;
1761 : out <= 12'b000000110100;
1762 : out <= 12'b000000110100;
1763 : out <= 12'b000000110100;
1764 : out <= 12'b000000110100;
1765 : out <= 12'b000000110011;
1766 : out <= 12'b000000110011;
1767 : out <= 12'b000000110011;
1768 : out <= 12'b000000110011;
1769 : out <= 12'b000000110011;
1770 : out <= 12'b000000110011;
1771 : out <= 12'b000000110011;
1772 : out <= 12'b000000110011;
1773 : out <= 12'b000000110011;
1774 : out <= 12'b000000110011;
1775 : out <= 12'b000000110011;
1776 : out <= 12'b000000110011;
1777 : out <= 12'b000000110011;
1778 : out <= 12'b000000110011;
1779 : out <= 12'b000000110011;
1780 : out <= 12'b000000110011;
1781 : out <= 12'b000000110011;
1782 : out <= 12'b000000110011;
1783 : out <= 12'b000000110011;
1784 : out <= 12'b000000110011;
1785 : out <= 12'b000000110011;
1786 : out <= 12'b000000110011;
1787 : out <= 12'b000000110011;
1788 : out <= 12'b000000110011;
1789 : out <= 12'b000000110011;
1790 : out <= 12'b000000110011;
1791 : out <= 12'b000000110011;
1792 : out <= 12'b000000110011;
1793 : out <= 12'b000000110011;
1794 : out <= 12'b000000110011;
1795 : out <= 12'b000000110011;
1796 : out <= 12'b000000110011;
1797 : out <= 12'b000000110011;
1798 : out <= 12'b000000110011;
1799 : out <= 12'b000000110011;
1800 : out <= 12'b000000110011;
1801 : out <= 12'b000000110011;
1802 : out <= 12'b000000110011;
1803 : out <= 12'b000000110011;
1804 : out <= 12'b000000110011;
1805 : out <= 12'b000000110011;
1806 : out <= 12'b000000110011;
1807 : out <= 12'b000000110011;
1808 : out <= 12'b000000110011;
1809 : out <= 12'b000000110011;
1810 : out <= 12'b000000110011;
1811 : out <= 12'b000000110011;
1812 : out <= 12'b000000110011;
1813 : out <= 12'b000000110011;
1814 : out <= 12'b000000110011;
1815 : out <= 12'b000000110011;
1816 : out <= 12'b000000110011;
1817 : out <= 12'b000000110011;
1818 : out <= 12'b000000110011;
1819 : out <= 12'b000000110010;
1820 : out <= 12'b000000110010;
1821 : out <= 12'b000000110010;
1822 : out <= 12'b000000110010;
1823 : out <= 12'b000000110010;
1824 : out <= 12'b000000110010;
1825 : out <= 12'b000000110010;
1826 : out <= 12'b000000110010;
1827 : out <= 12'b000000110010;
1828 : out <= 12'b000000110010;
1829 : out <= 12'b000000110010;
1830 : out <= 12'b000000110010;
1831 : out <= 12'b000000110010;
1832 : out <= 12'b000000110010;
1833 : out <= 12'b000000110010;
1834 : out <= 12'b000000110010;
1835 : out <= 12'b000000110010;
1836 : out <= 12'b000000110010;
1837 : out <= 12'b000000110010;
1838 : out <= 12'b000000110010;
1839 : out <= 12'b000000110010;
1840 : out <= 12'b000000110010;
1841 : out <= 12'b000000110010;
1842 : out <= 12'b000000110010;
1843 : out <= 12'b000000110010;
1844 : out <= 12'b000000110010;
1845 : out <= 12'b000000110010;
1846 : out <= 12'b000000110010;
1847 : out <= 12'b000000110010;
1848 : out <= 12'b000000110010;
1849 : out <= 12'b000000110010;
1850 : out <= 12'b000000110010;
1851 : out <= 12'b000000110010;
1852 : out <= 12'b000000110010;
1853 : out <= 12'b000000110010;
1854 : out <= 12'b000000110010;
1855 : out <= 12'b000000110010;
1856 : out <= 12'b000000110010;
1857 : out <= 12'b000000110010;
1858 : out <= 12'b000000110010;
1859 : out <= 12'b000000110010;
1860 : out <= 12'b000000110010;
1861 : out <= 12'b000000110010;
1862 : out <= 12'b000000110010;
1863 : out <= 12'b000000110010;
1864 : out <= 12'b000000110010;
1865 : out <= 12'b000000110010;
1866 : out <= 12'b000000110010;
1867 : out <= 12'b000000110010;
1868 : out <= 12'b000000110010;
1869 : out <= 12'b000000110010;
1870 : out <= 12'b000000110010;
1871 : out <= 12'b000000110010;
1872 : out <= 12'b000000110010;
1873 : out <= 12'b000000110010;
1874 : out <= 12'b000000110010;
1875 : out <= 12'b000000110010;
1876 : out <= 12'b000000110001;
1877 : out <= 12'b000000110001;
1878 : out <= 12'b000000110001;
1879 : out <= 12'b000000110001;
1880 : out <= 12'b000000110001;
1881 : out <= 12'b000000110001;
1882 : out <= 12'b000000110001;
1883 : out <= 12'b000000110001;
1884 : out <= 12'b000000110001;
1885 : out <= 12'b000000110001;
1886 : out <= 12'b000000110001;
1887 : out <= 12'b000000110001;
1888 : out <= 12'b000000110001;
1889 : out <= 12'b000000110001;
1890 : out <= 12'b000000110001;
1891 : out <= 12'b000000110001;
1892 : out <= 12'b000000110001;
1893 : out <= 12'b000000110001;
1894 : out <= 12'b000000110001;
1895 : out <= 12'b000000110001;
1896 : out <= 12'b000000110001;
1897 : out <= 12'b000000110001;
1898 : out <= 12'b000000110001;
1899 : out <= 12'b000000110001;
1900 : out <= 12'b000000110001;
1901 : out <= 12'b000000110001;
1902 : out <= 12'b000000110001;
1903 : out <= 12'b000000110001;
1904 : out <= 12'b000000110001;
1905 : out <= 12'b000000110001;
1906 : out <= 12'b000000110001;
1907 : out <= 12'b000000110001;
1908 : out <= 12'b000000110001;
1909 : out <= 12'b000000110001;
1910 : out <= 12'b000000110001;
1911 : out <= 12'b000000110001;
1912 : out <= 12'b000000110001;
1913 : out <= 12'b000000110001;
1914 : out <= 12'b000000110001;
1915 : out <= 12'b000000110001;
1916 : out <= 12'b000000110001;
1917 : out <= 12'b000000110001;
1918 : out <= 12'b000000110001;
1919 : out <= 12'b000000110001;
1920 : out <= 12'b000000110001;
1921 : out <= 12'b000000110001;
1922 : out <= 12'b000000110001;
1923 : out <= 12'b000000110001;
1924 : out <= 12'b000000110001;
1925 : out <= 12'b000000110001;
1926 : out <= 12'b000000110001;
1927 : out <= 12'b000000110001;
1928 : out <= 12'b000000110001;
1929 : out <= 12'b000000110001;
1930 : out <= 12'b000000110001;
1931 : out <= 12'b000000110001;
1932 : out <= 12'b000000110001;
1933 : out <= 12'b000000110001;
1934 : out <= 12'b000000110001;
1935 : out <= 12'b000000110001;
1936 : out <= 12'b000000110000;
1937 : out <= 12'b000000110000;
1938 : out <= 12'b000000110000;
1939 : out <= 12'b000000110000;
1940 : out <= 12'b000000110000;
1941 : out <= 12'b000000110000;
1942 : out <= 12'b000000110000;
1943 : out <= 12'b000000110000;
1944 : out <= 12'b000000110000;
1945 : out <= 12'b000000110000;
1946 : out <= 12'b000000110000;
1947 : out <= 12'b000000110000;
1948 : out <= 12'b000000110000;
1949 : out <= 12'b000000110000;
1950 : out <= 12'b000000110000;
1951 : out <= 12'b000000110000;
1952 : out <= 12'b000000110000;
1953 : out <= 12'b000000110000;
1954 : out <= 12'b000000110000;
1955 : out <= 12'b000000110000;
1956 : out <= 12'b000000110000;
1957 : out <= 12'b000000110000;
1958 : out <= 12'b000000110000;
1959 : out <= 12'b000000110000;
1960 : out <= 12'b000000110000;
1961 : out <= 12'b000000110000;
1962 : out <= 12'b000000110000;
1963 : out <= 12'b000000110000;
1964 : out <= 12'b000000110000;
1965 : out <= 12'b000000110000;
1966 : out <= 12'b000000110000;
1967 : out <= 12'b000000110000;
1968 : out <= 12'b000000110000;
1969 : out <= 12'b000000110000;
1970 : out <= 12'b000000110000;
1971 : out <= 12'b000000110000;
1972 : out <= 12'b000000110000;
1973 : out <= 12'b000000110000;
1974 : out <= 12'b000000110000;
1975 : out <= 12'b000000110000;
1976 : out <= 12'b000000110000;
1977 : out <= 12'b000000110000;
1978 : out <= 12'b000000110000;
1979 : out <= 12'b000000110000;
1980 : out <= 12'b000000110000;
1981 : out <= 12'b000000110000;
1982 : out <= 12'b000000110000;
1983 : out <= 12'b000000110000;
1984 : out <= 12'b000000110000;
1985 : out <= 12'b000000110000;
1986 : out <= 12'b000000110000;
1987 : out <= 12'b000000110000;
1988 : out <= 12'b000000110000;
1989 : out <= 12'b000000110000;
1990 : out <= 12'b000000110000;
1991 : out <= 12'b000000110000;
1992 : out <= 12'b000000110000;
1993 : out <= 12'b000000110000;
1994 : out <= 12'b000000110000;
1995 : out <= 12'b000000110000;
1996 : out <= 12'b000000110000;
1997 : out <= 12'b000000110000;
1998 : out <= 12'b000000110000;
1999 : out <= 12'b000000110000;
2000 : out <= 12'b000000110000;
	  default out<= 12'b000000000000;	
		
	  endcase
        
end 
 endmodule