module LEDLamp ( input clk,
	     input pulse,
	     output  LED);

COUNTER500 Counter00(clk,pulse,LED);

endmodule

module COUNTER500(input clk,      
                  input rstn,                
		  output reg allow);

 reg[10:0] out = 500 ;   

 always @ (posedge clk) begin  
    if ( rstn) begin 
      	out <= 0 ;
 	allow<=1;
	end	
    else if(out >= 500)
	allow <= 0;		  
    else  
      out <= out + 1 ;  
  end  

endmodule
