 
`timescale 1ms/100us 

module Test;

// ????? ??
reg clk ;
reg pulse ;
reg mute ;
reg start; // ????? ?? ?? ??? ?? ??? ???? ???? ???? ??? ?????? ???? ?????? ??? ???? ???? ???? ??? ???? ????? ??


// ??? ??? ????? ????? ??? ??? ??????
wire z ;       
wire[10:0] out;
wire[10:0] out1;
wire[11:0] out2;

// ????? ??
wire[6:0] seg0,seg1,seg2;
wire LED;
wire Speaker;

// ???? ????
always #0.5 clk = ~clk;

// ??? ??? ????? ???? ??? ???? ?? ??? ?

Pulse_finder PULSE_FINDER( clk,pulse,z); // ????? ?? ????? ???

LEDLamp LEDLAMP( clk,z,LED); // ?????? ?? ?? ??
Speaker_Controler SPEAKER_CONTROLER(mute,Speaker,clk,LED,start); // ?????? ??????

counter COUNTER( clk, z , out); // ??????? ?????
Register REGISTER( out,clk,z,out1); // ?????? ????? ????? ???
Rom ROM(out2,out1,clk); // eprom
segment7 SEG1(out2[3:0],seg0),SEG2(out2[7:4],seg1),SEG3(out2[11:8],seg2); // ??? ????? ??



 //  ??? ????
  initial begin  

    	clk <= 0; 
	pulse <=0; 
	mute <=0;
	start <=0;

	#(10) start = ~start;
	#(10) start = ~start;
	#(5)  pulse = ~pulse;
	#(10) pulse = ~pulse;
	#(10) mute = ~mute;
        #(10) mute = ~mute;
	#(400) mute = ~mute;
	#(10) mute = ~mute;
	#(427) pulse = ~pulse;
	#(10) pulse = ~pulse;
	#(987)pulse = ~pulse;
	#(10)pulse = ~pulse;
  end  
endmodule
